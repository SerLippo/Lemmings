`ifndef LEMMINGS_SEQUENCES_SVH
`define LEMMINGS_SEQUENCES_SVH

// elem seq
`include "lemmings_master_sequence.sv"

// virt seq
`include "lemmings_base_virtual_sequence.sv"
`include "lemmings_full_random_virt_seq.sv"
`include "lemmings_left_splat_virt_seq.sv"
`include "lemmings_right_splat_virt_seq.sv"

`endif
`ifndef LEMMINGS_DEFINE_SV
`define LEMMINGS_DEFINE_SV

typedef enum {LEFT, RIGHT, DIG_L, DIG_R, FALL_L, FALL_R, SPLAT} state_t;

`endif
`ifndef LEMMINGS_TESTS_SVH
`define LEMMINGS_TESTS_SVH

`include "lemmings_base_test.sv"
`include "lemmings_full_random_test.sv"
`include "lemmings_left_splat_test.sv"
`include "lemmings_right_splat_test.sv"

`endif